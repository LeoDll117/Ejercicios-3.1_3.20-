----------------------------------------------------------------------------------
--Ejercicio 3.5
--Leonardo Peralta 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;



entity Ejer35 is
    Port ( clk : in  STD_LOGIC;
           Q : inout  STD_LOGIC_VECTOR (5 downto 0);
           ns : out  STD_LOGIC_VECTOR (2 downto 0);
           eo : out  STD_LOGIC_VECTOR (2 downto 0);
           m : in  STD_LOGIC);
end Ejer35;

architecture Behavioral of Ejer35 is

begin


end Behavioral;

